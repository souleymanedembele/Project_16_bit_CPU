/**
 * File              : Processor.sv
 */

